b0VIM 8.0      �x�_J  �)  jetbot                                  jetson-4-3                              ~jetbot/catkin_ws/src/raspimouse_navigation_3/param/local_costmap_params.yaml                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                utf-8U3210    #"! U                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 tp                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        ad  �  �            �  �  �  �  �  s  e  R  >  '    �  �  �  �  D  �  �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  # - {name: obstacle_layer,       type: "costmap_2d::ObstacleLayer"}   # - {name: static_map,       type: "costmap_2d::StaticLayer"}   # - {name: inflation_layer,      type: "costmap_2d::InflationLayer"}   #plugins:    inflation_radius: 0.1   cost_scaling_factor: 0.5   transform_tolerance: 10.0   rolling_window: true   static_map: false   resolution: 0.01   height: 4.0   width: 4.0   publish_frequency: 10.0 #2.0   update_frequency: 10.0 #5.0   robot_base_frame: base_link   global_frame: odom local_costmap:  